module quick_rs232 #(
)
()

endmodule
